`timescale 1ns / 1ps
`include "processor_ci_defines.vh"
// `define ENABLE_SECOND_MEMORY 1

module processorci_top (
    `ifdef DIFERENCIAL_CLK
    input  logic clk_ref_p,
    input  logic clk_ref_n,
    `else
    input  logic clk,
    `endif

    input  logic rst,

    // UART pins
    input  logic rx,
    output logic tx
    `ifndef DIFERENCIAL_CLK
    ,

    // SPI pins
    input  logic sck,
    input  logic cs,
    input  logic mosi,
    output logic miso,

    //SPI control pins
    input  logic rw,
    output logic intr
    `endif
);

logic clk_o, rst_n;
logic clk_core, rst_core;


// Fios do barramento entre Controller e Processor
logic        core_cyc;
logic        core_stb;
logic        core_we;
logic [31:0] core_addr;
logic [31:0] core_data_out;
logic [31:0] core_data_in;
logic        core_ack;

`ifdef ENABLE_SECOND_MEMORY
logic        data_mem_cyc;
logic        data_mem_stb;
logic        data_mem_we;
logic [31:0] data_mem_addr;
logic [31:0] data_mem_data_out;
logic [31:0] data_mem_data_in;
logic        data_mem_ack;
`endif


Controller #(
    .CLK_FREQ           (`CLOCK_FREQ),
    .BIT_RATE           (`BIT_RATE),
    .PAYLOAD_BITS       (`PAYLOAD_BITS),
    .BUFFER_SIZE        (`BUFFER_SIZE),
    .PULSE_CONTROL_BITS (`PULSE_CONTROL_BITS),
    .BUS_WIDTH          (`BUS_WIDTH),
    .WORD_SIZE_BY       (`WORD_SIZE_BY),
    .ID                 (`ID),
    .RESET_CLK_CYCLES   (`RESET_CLK_CYCLES),
    .MEMORY_FILE        (`MEMORY_FILE),
    .MEMORY_SIZE        (`MEMORY_SIZE)
) u_Controller (
    `ifdef HIGH_CLK
    .clk                (clk_o),
    `else
    .clk                (clk),
    `endif

    .rst_n              (rst_n),
    
    // SPI signals
    .sck_i              (sck),
    .cs_i               (cs),
    .mosi_i             (mosi),
    .miso_o             (miso),
    
    // SPI callback signals
    .rw_i               (rw),
    .intr_o             (intr),
    
    // UART signals
    .rx                 (rx),
    .tx                 (tx),
    
    // Clock, reset, and bus signals
    .clk_core_o         (clk_core),
    .rst_core_o         (rst_core),
    
    // Barramento padrão (Wishbone)
    .core_cyc_i         (core_cyc),
    .core_stb_i         (core_stb),
    .core_we_i          (core_we),
    .core_addr_i        (core_addr),
    .core_data_i        (core_data_out),
    .core_data_o        (core_data_in),
    .core_ack_o         (core_ack)

    `ifdef ENABLE_SECOND_MEMORY
    ,
    .data_mem_cyc_i     (data_mem_cyc),
    .data_mem_stb_i     (data_mem_stb),
    .data_mem_we_i      (data_mem_we),
    .data_mem_addr_i    (data_mem_addr),
    .data_mem_data_i    (data_mem_data_out),
    .data_mem_data_o    (data_mem_data_in),
    .data_mem_ack_o     (data_mem_ack)
    `endif
);

// Core space

neorv32_cpu #(
  // General
  .HART_ID              (0),
  .BOOT_ADDR            (32'h00000000),
  .DEBUG_PARK_ADDR      (32'h00000000),
  .DEBUG_EXC_ADDR       (32'h00000000),
  .ICC_EN               (1'b1),

  // RISC-V ISA Extensions
  .RISCV_ISA_C          (1'b1),
  .RISCV_ISA_E          (1'b1),
  .RISCV_ISA_M          (1'b1),
  .RISCV_ISA_U          (1'b1),
  .RISCV_ISA_Zaamo      (1'b1),
  .RISCV_ISA_Zalrsc     (1'b1),
  .RISCV_ISA_Zba        (1'b1),
  .RISCV_ISA_Zbb        (1'b1),
  .RISCV_ISA_Zbkb       (1'b1),
  .RISCV_ISA_Zbkc       (1'b1),
  .RISCV_ISA_Zbkx       (1'b1),
  .RISCV_ISA_Zbs        (1'b1),
  .RISCV_ISA_Zfinx      (1'b1),
  .RISCV_ISA_Zicntr     (1'b1),
  .RISCV_ISA_Zicond     (1'b1),
  .RISCV_ISA_Zihpm      (1'b1),
  .RISCV_ISA_Zknd       (1'b1),
  .RISCV_ISA_Zkne       (1'b1),
  .RISCV_ISA_Zknh       (1'b1),
  .RISCV_ISA_Zksed      (1'b1),
  .RISCV_ISA_Zksh       (1'b1),
  .RISCV_ISA_Zmmul      (1'b1),
  .RISCV_ISA_Zxcfu      (1'b1),
  .RISCV_ISA_Sdext      (1'b1),
  .RISCV_ISA_Sdtrig     (1'b1),
  .RISCV_ISA_Smpmp      (1'b1),

  // Tuning Options
  .CPU_FAST_MUL_EN      (1'b1),
  .CPU_FAST_SHIFT_EN    (1'b1),
  .CPU_RF_HW_RST_EN     (1'b1),

  // Physical Memory Protection (PMP)
  .PMP_NUM_REGIONS      (16),
  .PMP_MIN_GRANULARITY  (64),
  .PMP_TOR_MODE_EN      (1'b1),
  .PMP_NAP_MODE_EN      (1'b1),

  // Hardware Performance Monitors (HPM)
  .HPM_NUM_CNTS         (13),
  .HPM_CNT_WIDTH        (64)
) u_neorv32_cpu (
  // Global control
  .clk_i                (clk_core),
  .rstn_i               (rst_core),

  // Interrupts
  .msi_i                (),
  .mei_i                (),
  .mti_i                (),
  .firq_i               (),
  .dbi_i                (),

  // Inter-core communication links
  .icc_tx_o             (),
  .icc_rx_i             (),

  // Instruction bus interface
  .ibus_req_o           (),
  .ibus_rsp_i           (),

  // Data bus interface
  .dbus_req_o           (),
  .dbus_rsp_i           (),

  // Memory synchronization
  .mem_sync_i           ()
);

// Clock inflaestructure

initial begin
    clk_o = 1'b0; // 50mhz or 100mhz
end

`ifdef DIFERENCIAL_CLK
logic clk_ref; // Sinal de clock single-ended

// Differential clock input
IBUFDS #(
    .DIFF_TERM    ("FALSE"), // Enable or disable differential terminator
    .IBUF_LOW_PWR ("TRUE"),  // Enable low power mode
    .IOSTANDARD   ("DIFF_SSTL15")
) ibufds_inst (
    .O  (clk_ref),   // Clock single-ended output
    .I  (clk_ref_p), // Differential input positive
    .IB (clk_ref_n)  // Differential input negative
);


always_ff @(posedge clk_ref) begin
    clk_o <= ~clk_o;
end
`else
always_ff @(posedge clk) begin
    clk_o <= ~clk_o;
end
`endif


// Reset Inflaestructure


ResetBootSystem #(
    .CYCLES(20)
) ResetBootSystem(
    `ifdef HIGH_CLK
    .clk     (clk_o),
    `else
    .clk     (clk),
    `endif
    
    .rst_n_o (rst_n)
);
    
endmodule
